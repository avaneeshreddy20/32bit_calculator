library ieee;
use ieee.std_logic_1164.all;
entity ff is
  port ( a : in std_logic;
         load,clear,clock : in std_logic;
         z : out std_logic );
end ff;
architecture behavioural of ff is
begin
  process(clear,clock)
    begin
  if (clear = '1') then
    z <= '0' ;
  elsif (rising_edge(clock)) then
   if ( load = '1' ) then 
  z <= a;
end if;
  end if;
  end process;
end behavioural;
