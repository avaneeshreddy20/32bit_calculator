library ieee;
use ieee.std_logic_1164.all;
entity divider is
  port ( a  : in std_logic_vector( 15 downto 0);
         c  : out std_logic_vector(15 downto 0));
end divider;

architecture structural of divider is
begin
  c <= "00" & a(15 downto 2);
end structural;